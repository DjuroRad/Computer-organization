`define CLOCK 4
`define DELAY 1250
module alu_32bit_with_mult_testbench();


	//module mult_64bit(product, a, b, clk);

	reg [31:0] a, b;
	reg clk;
	reg [2:0]alu_op;
	wire [31:0] res;

	alu_32bit_with_mult alumult32(res, alu_op, a, b, clk);
	
	initial begin
	clk = 1'b0;
	//mult
	alu_op = 3'b011; a =32'b0000_0000_0000_0000_0000_0000_0000_1111; b = 32'b0000_0000_0000_0000_0000_0000_0000_0011;
	#`DELAY;
	//add
	alu_op = 3'b000; a =32'b0000_0000_0000_0000_0000_0000_0000_1101; b = 32'b0000_0000_0000_0000_0000_0000_0000_1100;
	#`DELAY;
	//xor
	alu_op = 3'b001; a =32'b0000_0010_0000_0000_0000_0000_0000_1101; b = 32'b0000_0010_0000_0000_0000_0000_0000_1100;
	#`DELAY;
	//sub
	alu_op = 3'b010; a =32'b0000_0000_0000_0000_0000_0000_0000_1101; b = 32'b0000_0000_0000_0000_0000_0000_0000_0111;
	#`DELAY;
	//sub
	alu_op = 3'b010; a =32'b1000_0000_0000_0000_0000_0000_0000_1101; b = 32'b1000_0000_0000_0000_0000_0000_0000_1111;
	#`DELAY;
	//slt
	alu_op = 3'b100; a =32'b0000_0010_0000_0000_0000_0000_0000_1101; b = 32'b0000_0010_0000_0000_0000_0000_0000_1100;
	#`DELAY;
	//slt
	alu_op = 3'b100; a =32'b0000_0010_0000_0000_0000_0000_0000_1101; b = 32'b0010_0010_0000_0000_0000_0000_0000_1100;
	#`DELAY;
	//nor
	alu_op = 3'b101; a =32'b0000_0010_0000_0000_0000_0000_0000_1101; b = 32'b0000_0010_0000_0000_0000_0000_0000_1100;
	#`DELAY;
	//and
	alu_op = 3'b110; a =32'b0000_0010_0000_0000_0000_0000_0000_1101; b = 32'b0000_0010_0000_0000_0000_0000_0000_1100;
	#`DELAY;
	//or
	alu_op = 3'b111; a =32'b0000_0010_0000_0000_0000_0000_0000_1101; b = 32'b0000_0010_0000_0000_0000_0000_0000_1100;
	#`DELAY;
	#2000 $finish;
	end
	
	//define clock cycle
	always
		begin
			#4 clk = ~clk;
		end
		
	initial begin
	$monitor("time=%2d, res=%32b, a=%32b, b=%32b"
	          ,$time, res, a, b);
	end
	
	

endmodule