module control_unit_multiplier(next_state, state, i_eq_0, p_lsb, a_sel);
input [2:0]next_state, state;
input i_eq_0, p_lsb, a_sel;

//not(a_not, a);
//not(b_not, b);

//and( a_b_not, a, b_not );
//and( a_not_b, a_not, b);

//or( res, a_b_not, a_not_b );

endmodule