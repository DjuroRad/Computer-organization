library verilog;
use verilog.vl_types.all;
entity \_xor\ is
    port(
        res             : out    vl_logic;
        a               : in     vl_logic;
        b               : in     vl_logic
    );
end \_xor\;
