`define DELAY 20
module alu_32bit_testbench();
	
	reg [31:0] a, b;
	reg [2:0] alu_op;
	wire [31:0]res;
	wire zero;
	//module module alu_32bit(res, alu_op, a, b);
	alu_32bit alu32bit(res, alu_op , a, b, zero);
	
	initial begin
	//add
	alu_op = 3'b000; a =32'b0000_0000_0000_0000_0000_0000_0000_1101; b = 32'b0000_0000_0000_0000_0000_0000_0000_1100;
	#`DELAY;
	//xor
	alu_op = 3'b001; a =32'b0000_0010_0000_0000_0000_0000_0000_1101; b = 32'b0000_0010_0000_0000_0000_0000_0000_1100;
	#`DELAY;
	//sub
	alu_op = 3'b010; a =32'b0000_0000_0000_0000_0000_0000_0000_1101; b = 32'b0000_0000_0000_0000_0000_0000_0000_0111;
	#`DELAY;
	//sub
	alu_op = 3'b010; a =32'b1000_0000_0000_0000_0000_0000_0000_1101; b = 32'b1000_0000_0000_0000_0000_0000_0000_1111;
	#`DELAY;
	//sub
	alu_op = 3'b010; a =32'b1000_0000_0000_0000_0000_0000_0000_1101; b = 32'b1000_0000_0000_0000_0000_0000_0000_1101;
	#`DELAY
	//mult
	alu_op = 3'b011; a =32'b0000_0000_0000_0000_0000_0000_0000_1101; b = 32'b0000_0000_0000_0000_0000_0000_0000_1100;
	#`DELAY;
	//slt
	alu_op = 3'b100; a =32'b0000_0010_0000_0000_0000_0000_0000_1101; b = 32'b0000_0010_0000_0000_0000_0000_0000_1100;
	#`DELAY;
	//slt
	alu_op = 3'b100; a =32'b0000_0010_0000_0000_0000_0000_0000_1101; b = 32'b0010_0010_0000_0000_0000_0000_0000_1100;
	#`DELAY;
	//nor
	alu_op = 3'b101; a =32'b0000_0010_0000_0000_0000_0000_0000_1101; b = 32'b0000_0010_0000_0000_0000_0000_0000_1100;
	#`DELAY;
	//and
	alu_op = 3'b110; a =32'b0000_0010_0000_0000_0000_0000_0000_1101; b = 32'b0000_0010_0000_0000_0000_0000_0000_1100;
	#`DELAY;
	//or
	alu_op = 3'b111; a =32'b0000_0010_0000_0000_0000_0000_0000_1101; b = 32'b0000_0010_0000_0000_0000_0000_0000_1100;
	#`DELAY;
	end
	initial begin
	$monitor("time=%2d,a=%32b,b=%32b alu_op2=%1b,alu_op1=%1b,alu_op0=%1b,res=%32b"
	          ,$time, a, b, alu_op[2], alu_op[1], alu_op[0], res);
	end
endmodule